`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:07:18 04/15/2019 
// Design Name: 
// Module Name:    fixedfloat 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fixedfloat(
    input clk,
    input rst,
    input targetnumber,
    input fixpointpos,
    input opcode,
    output result
    );


endmodule
