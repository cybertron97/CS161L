`timescale 1ns / 1ps

module myalutb;

	parameter NUMBITS = 8 ;

	// Inputs
	reg clk ;
	reg reset ; 
	reg [NUMBITS-1:0] A;
	reg [NUMBITS-1:0] B;
	reg [2:0] opcode;

	// Outputs
	
	wire [NUMBITS-1:0] result;
	reg [NUMBITS-1:0] R ;
	wire carryout;
	wire overflow;
	wire zero;

   // -------------------------------------------------------
	// Instantiate the Unit Under Test (UUT)
	// -------------------------------------------------------
	
	my_alu #(NUMBITS) uut (
	   .clk(clk),
		.reset(reset) ,  
		.A(A), 
		.B(B), 
		.opcode(opcode), 
		.result(result), 
		.carryout(carryout), 
		.overflow(overflow), 
		.zero(zero)
	);

  	initial begin 
	
	 clk = 0 ; reset = 1 ; #50 ; 
	 clk = 1 ; reset = 1 ; #50 ; 
	 clk = 0 ; reset = 0 ; #50 ; 
	 clk = 1 ; reset = 0 ; #50 ; 
		 
	 forever begin 
		clk = ~clk; #50 ; 
	 end 
	 
	end 
	
	initial begin
		
		// ---------------------------------------------
		// Testing unsigned additions 
		// --------------------------------------------- 
		opcode = 3'b000 ; 
		A = 8'hFF ;
   	B = 8'h01 ;
		R = 8'h00 ; 
		
	    #100 ; // Wait 
     
		$display("TC11 Unsigned Add ");
		if (R != result) $display  ("Result is wrong");
		if (zero != 1'b1) $display ("Zero  is wrong");
		if (carryout != 1'b1) $display ("Carryout is wrong");
		
		A = 8'h01 ;
   	B = 8'h00 ;
		R = 8'h01 ; 
		
	    #100 ; // Wait 
     
		$display("TC12 Unsigned Add ");
		if (R != result) $display  ("Result is wrong");
		if (zero != 1'b0) $display ("Zero  is wrong");
		if (carryout != 1'b0) $display ("Carryout is wrong");
		
		A = 8'hff ;
   	B = 8'h01 ;
		R = 8'h00 ; 
		
	    #100 ; // Wait 
     
		$display("TC13 Unsigned Add ");
		if (R != result) $display  ("Result is wrong");
		if (zero != 1'b1) $display ("Zero  is wrong");
		if (carryout != 1'b1) $display ("Carryout is wrong");
		
		A = 8'h0f ;
   	B = 8'hf0 ;
		R = 8'hff ; 
		
	    #100 ; // Wait 
     
		$display("TC14 Unsigned Add ");
		if (R != result) $display  ("Result is wrong");
		if (zero != 1'b0) $display ("Zero  is wrong");
		if (carryout != 1'b0) $display ("Carryout is wrong");
		
		A = 8'h0f ;
   	B = 8'h0f ;
		R = 8'h1e ; 
		
	    #100 ; // Wait 
     
		$display("TC15 Unsigned Add ");
		if (R != result) $display  ("Result is wrong");
		if (zero != 1'b0) $display ("Zero  is wrong");
		if (carryout != 1'b0) $display ("Carryout is wrong");
		
		
		
		
		// ---------------------------------------------
		// Testing unsigned subs 
		// --------------------------------------------- 

       opcode= 3'b010; 
		 A = 8'h00 ;
   	 B = 8'h00 ;
		 R = 8'h00 ; 
		
	    #100 ; // Wait 
     
		$display("TC16 Unsigned subs ");
		if (R != result) $display  ("Result is wrong");
		if (zero != 1'b1) $display ("Zero  is wrong");
		if (carryout != 1'b0) $display ("Carryout is wrong");
		
		 A = 8'hff ;
   	 B = 8'hff ;
		 R = 8'h00 ; 
		
	    #100 ; // Wait 
     
		$display("TC17 Unsigned subs ");
		if (R != result) $display  ("Result is wrong");
		if (zero != 1'b1) $display ("Zero  is wrong");
		if (carryout != 1'b0) $display ("Carryout is wrong");
		
		 A = 8'h1f ;
   	 B = 8'h0f ;
		 R = 8'h10 ; 
		
	    #100 ; // Wait 
     
		$display("TC18 Unsigned subs ");
		if (R != result) $display  ("Result is wrong");
		if (zero != 1'b0) $display ("Zero  is wrong");
		if (carryout != 1'b0) $display ("Carryout is wrong");
		
		 A = 8'h0A ;
   	 B = 8'h01 ;
		 R = 8'h09 ; 
		
	    #100 ; // Wait 
     
		$display("TC19 Unsigned subs ");
		if (R != result) $display  ("Result is wrong");
		if (zero != 1'b0) $display ("Zero  is wrong");
		if (carryout != 1'b0) $display ("Carryout is wrong");
		
		// ---------------------------------------------
		// Testing signed adds 
		// --------------------------------------------- 
		opcode = 3'b001; 
		
		A=8'h0A;
		B=8'h01;
		R=8'h0B;
		
		#100; 
		$display("TC20 signed adds ");
		if (R != result) $display  ("Result is wrong");
		if (zero != 1'b0) $display ("Zero  is wrong");
		if (carryout != 1'b0) $display ("Carryout is wrong");
		
		A=8'hAE;
		B=8'h01;
		R=8'hAF;
		
		#100; 
		$display("TC21 signed adds ");
		if (R != result) $display  ("Result is wrong");
		if (zero != 1'b0) $display ("Zero  is wrong");
		if (carryout != 1'b0) $display ("Carryout is wrong");
		
		A=8'hAE;
		B=$signed(~({8'hAE}))+$signed(2'b01);
		R=8'h00;
		
		#100; 
		$display("TC22 signed adds ");
		if (R != result) $display  ("Result is wrong");
		if (zero != 1'b1) $display ("Zero  is wrong");
		if (carryout != 1'b0) $display ("Carryout is wrong");
		
		// ---------------------------------------------
		// Testing signed subs 
		// --------------------------------------------- 
		
		// ---------------------------------------------
		// Testing ANDS 
		// --------------------------------------------- 
		
		// ----------------------------------------
		// ORs 
		// ---------------------------------------- 
		
		// ----------------------------------------
		// XORs 
		// ---------------------------------------- 

		// ----------------------------------------
		// Div 2 
		// ----------------------------------------
	end
      
endmodule
